module _not(output y, input a);    
    not(y, a);
endmodule