module _not(output y, input a);
    nand(y, a, a);
endmodule