module _and(output y, input a, b);    
    and(y, a, b);
endmodule